library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

--TODO THIS IS JUST A NORMAL REGISTER RIGHT NOW (NEED TO ADAPT FOR PIPELINE)
entity EXMEM is
    Port (
        clk        : in  STD_LOGIC;
        i_RST      : in  STD_LOGIC;
        reg_write  : in  STD_LOGIC;
        write_alu_data : in  STD_LOGIC_VECTOR (31 downto 0);
        write_aluSrc_data : in  STD_LOGIC_VECTOR (31 downto 0); --Not sure if this is what the input is actually coming from need to double check
        write_wrMuxO_data : in STD_LOGIC_VECTOR(4 downto 0);
        write_nextAddr_data : in STD_LOGIC_VECTOR(31 downto 0);
        write_reg2out_data : in STD_LOGIC_VECTOR(31 downto 0);
        write_currentInstruction_data : in STD_LOGIC_VECTOR(31 downto 0);
        read_alu_data : out STD_LOGIC_VECTOR (31 downto 0);
        read_aluSrc_data : out STD_LOGIC_VECTOR (31 downto 0);
        read_wrMuxO_data : out STD_LOGIC_VECTOR(31 downto 0);
        read_nextAddr_data : out STD_LOGIC_VECTOR(31 downto 0);
        read_reg2out_data : out STD_LOGIC_VECTOR(31 downto 0);
        read_currentInstruction_data : out STD_LOGIC_VECTOR(31 downto 0);
        halt : in std_logic
    );
end EXMEM;


architecture Behavioral of EXMEM is
    type reg_array is array (0 to 31) of STD_LOGIC_VECTOR (31 downto 0);
    signal registers : reg_array := (others => (others => '0'));
    signal write_alu_reg : std_logic_vector(4 downto 0) := "00001";
    signal write_aluSrc_reg : std_logic_vector(4 downto 0) := "00010";
    signal write_wrMuxO_reg : std_logic_vector(4 downto 0) := "00011";
    signal write_nextAddr_reg : STD_LOGIC_VECTOR(4 downto 0) := "00100";
    signal write_reg2out_reg : STD_LOGIC_VECTOR(4 downto 0) := "00110";
    signal write_currentInstruction_reg : STD_LOGIC_VECTOR(4 downto 0) := "00111";
    signal write_aluBmux_reg : STD_LOGIC_VECTOR(4 downto 0) := "01111";
begin
    process(clk)
    begin
        if rising_edge(clk) then
            if i_RST = '1' then
                for i in 1 to 31 loop
                    registers(i) <= (others => '0');
                end loop;
            elsif (reg_write = '1' and halt = '0')  then                
                registers(to_integer(unsigned(write_alu_reg))) <= write_alu_data;
                registers(to_integer(unsigned(write_aluSrc_reg))) <= write_aluSrc_data;
                registers(to_integer(unsigned(write_wrMuxO_reg))) <= "000000000000000000000000000" & write_wrMuxO_data;
                registers(to_integer(unsigned(write_nextAddr_reg))) <= write_nextAddr_data;
                registers(to_integer(unsigned(write_reg2out_reg))) <= write_reg2out_data;
                registers(to_integer(unsigned(write_currentInstruction_reg))) <= write_currentInstruction_data;
            end if;
        end if;
    end process;
    read_alu_data <= registers(to_integer(unsigned(write_alu_reg)));
    read_aluSrc_data <= registers(to_integer(unsigned(write_aluSrc_reg)));
    read_wrMuxO_data <= registers(to_integer(unsigned(write_wrMuxO_reg)));
    read_nextAddr_data <= registers(to_integer(unsigned(write_nextAddr_reg)));
    read_reg2out_data <= registers(to_integer(unsigned(write_reg2out_reg)));
    read_currentInstruction_data <= registers(to_integer(unsigned(write_currentInstruction_reg)));
end Behavioral;

