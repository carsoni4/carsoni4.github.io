
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity pc_dff is

  port(
       i_CLK        : in std_logic;     -- Clock input
       i_RST        : in std_logic;     -- Reset input
       i_D          : in std_logic;     -- Data value input
       o_Q          : out std_logic;   -- Data value output
       i_RST_Data   : in std_logic;    -- Data input so we can initialize on rst
       halt  	    : in std_logic
       );   
end pc_dff;

architecture mixed of pc_dff is

  signal s_Q    : std_logic;    -- Output of the FF


begin

  -- The output of the FF is fixed to s_Q
  o_Q <= s_Q;

  
  --no more WE since its pc


  -- This process handles the asyncrhonous reset and
  -- synchronous write. We want to be able to reset 
  -- our processor's registers so that we minimize
  -- glitchy behavior on startup.
  process (i_CLK, i_RST)
  begin
    if (i_RST = '1') then
      s_Q <= i_RST_Data; -- Use "(others => '0')" for N-bit values
    elsif (rising_edge(i_CLK)) then
    	if halt = '0' then
      s_Q <= i_D; --since no WE doesnt matter
    	end if;
    end if;

  end process;
  
end mixed;
